module decoder4x16 // 4 x 16 decoder
(
	input [3:0] in,
	output [15:0] out
);
reg [15:0] r_o;
assign out = r_o;
always@* begin
	case(in)
		4'b0000: r_o <= 16'b0000000000000001;
		4'b0001: r_o <= 16'b0000000000000010;
		4'b0010: r_o <= 16'b0000000000000100;
		4'b0011: r_o <= 16'b0000000000001000;
		4'b0100: r_o <= 16'b0000000000010000;
		4'b0101: r_o <= 16'b0000000000100000;
		4'b0110: r_o <= 16'b0000000001000000;
		4'b0111: r_o <= 16'b0000000010000000;
		4'b1000: r_o <= 16'b0000000100000000;
		4'b1001: r_o <= 16'b0000001000000000;
		4'b1010: r_o <= 16'b0000010000000000;
		4'b1011: r_o <= 16'b0000100000000000;
		4'b1100: r_o <= 16'b0001000000000000;
		4'b1101: r_o <= 16'b0010000000000000;
		4'b1110: r_o <= 16'b0100000000000000;
		4'b1111: r_o <= 16'b1000000000000000;
	endcase
end
endmodule